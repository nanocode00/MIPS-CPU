module hello;
    initial begin
        $display("Hello, Verilog!");
        $finish;
    end
endmodule
