module Opcode_Decoder(
    input [5:0] op,
    output MemRead,
    output MemWrite,
    output ALUSrc,
    output Jump,
    output MemtoReg,
    output Branch,
    output RegDst,
    output RegWrite,
    output BneBeq,
    output IsJAL,
    output ZeroExtend
);

    wire RTYPE, J, JAL, BEQ, BNE, ADDI, ADDIU, SLTI, ANDI, ORI, XORI, COP0, LW, SW;

    assign RTYPE = op == 6'b000000;
    assign J     = op == 6'b000010;
    assign JAL   = op == 6'b000011;
    assign BEQ   = op == 6'b000100;
    assign BNE   = op == 6'b000101;
    assign ADDI  = op == 6'b001000;
    assign ADDIU = op == 6'b001001;
    assign SLTI  = op == 6'b001010;
    assign ANDI  = op == 6'b001100;
    assign ORI   = op == 6'b001101;
    assign XORI  = op == 6'b001110;
    assign COP0  = op == 6'b010000;
    assign LW    = op == 6'b100011;
    assign SW    = op == 6'b101011;

    assign MemRead    = LW;
    assign MemWrite   = SW;
    assign ALUSrc     = LW || SW || ANDI || ORI || SLTI || ADDIU || ADDI;
    assign Jump       = J || JAL;
    assign MemtoReg   = LW;
    assign Branch     = BEQ || BNE;
    assign RegDst     = RTYPE;
    assign RegWrite   = RTYPE || LW || ANDI || ORI || SLTI || ADDIU || ADDI || JAL || COP0;
    assign BneBeq     = BNE;
    assign IsJAL      = JAL;
    assign ZeroExtend = ANDI || ORI || XORI;

endmodule
